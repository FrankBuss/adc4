library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

entity crc8 is
	port (
		iCLK : in std_logic;

		init : in std_logic;
		update : in std_logic;
		data : in unsigned(7 downto 0);
		checksum : out unsigned(7 downto 0)
	);
end crc8;

architecture Behavior of crc8 is

	signal i_checksum : unsigned(7 downto 0);
	signal load_table : std_logic;

begin

	process (iCLK)
	begin
		if rising_edge(iCLK) then
			load_table <= '0';
			if load_table = '1' then
				case i_checksum is
					when x"00" => i_checksum <= x"00";
					when x"01" => i_checksum <= x"07";
					when x"02" => i_checksum <= x"0e";
					when x"03" => i_checksum <= x"09";
					when x"04" => i_checksum <= x"1c";
					when x"05" => i_checksum <= x"1b";
					when x"06" => i_checksum <= x"12";
					when x"07" => i_checksum <= x"15";
					when x"08" => i_checksum <= x"38";
					when x"09" => i_checksum <= x"3f";
					when x"0a" => i_checksum <= x"36";
					when x"0b" => i_checksum <= x"31";
					when x"0c" => i_checksum <= x"24";
					when x"0d" => i_checksum <= x"23";
					when x"0e" => i_checksum <= x"2a";
					when x"0f" => i_checksum <= x"2d";
					when x"10" => i_checksum <= x"70";
					when x"11" => i_checksum <= x"77";
					when x"12" => i_checksum <= x"7e";
					when x"13" => i_checksum <= x"79";
					when x"14" => i_checksum <= x"6c";
					when x"15" => i_checksum <= x"6b";
					when x"16" => i_checksum <= x"62";
					when x"17" => i_checksum <= x"65";
					when x"18" => i_checksum <= x"48";
					when x"19" => i_checksum <= x"4f";
					when x"1a" => i_checksum <= x"46";
					when x"1b" => i_checksum <= x"41";
					when x"1c" => i_checksum <= x"54";
					when x"1d" => i_checksum <= x"53";
					when x"1e" => i_checksum <= x"5a";
					when x"1f" => i_checksum <= x"5d";
					when x"20" => i_checksum <= x"e0";
					when x"21" => i_checksum <= x"e7";
					when x"22" => i_checksum <= x"ee";
					when x"23" => i_checksum <= x"e9";
					when x"24" => i_checksum <= x"fc";
					when x"25" => i_checksum <= x"fb";
					when x"26" => i_checksum <= x"f2";
					when x"27" => i_checksum <= x"f5";
					when x"28" => i_checksum <= x"d8";
					when x"29" => i_checksum <= x"df";
					when x"2a" => i_checksum <= x"d6";
					when x"2b" => i_checksum <= x"d1";
					when x"2c" => i_checksum <= x"c4";
					when x"2d" => i_checksum <= x"c3";
					when x"2e" => i_checksum <= x"ca";
					when x"2f" => i_checksum <= x"cd";
					when x"30" => i_checksum <= x"90";
					when x"31" => i_checksum <= x"97";
					when x"32" => i_checksum <= x"9e";
					when x"33" => i_checksum <= x"99";
					when x"34" => i_checksum <= x"8c";
					when x"35" => i_checksum <= x"8b";
					when x"36" => i_checksum <= x"82";
					when x"37" => i_checksum <= x"85";
					when x"38" => i_checksum <= x"a8";
					when x"39" => i_checksum <= x"af";
					when x"3a" => i_checksum <= x"a6";
					when x"3b" => i_checksum <= x"a1";
					when x"3c" => i_checksum <= x"b4";
					when x"3d" => i_checksum <= x"b3";
					when x"3e" => i_checksum <= x"ba";
					when x"3f" => i_checksum <= x"bd";
					when x"40" => i_checksum <= x"c7";
					when x"41" => i_checksum <= x"c0";
					when x"42" => i_checksum <= x"c9";
					when x"43" => i_checksum <= x"ce";
					when x"44" => i_checksum <= x"db";
					when x"45" => i_checksum <= x"dc";
					when x"46" => i_checksum <= x"d5";
					when x"47" => i_checksum <= x"d2";
					when x"48" => i_checksum <= x"ff";
					when x"49" => i_checksum <= x"f8";
					when x"4a" => i_checksum <= x"f1";
					when x"4b" => i_checksum <= x"f6";
					when x"4c" => i_checksum <= x"e3";
					when x"4d" => i_checksum <= x"e4";
					when x"4e" => i_checksum <= x"ed";
					when x"4f" => i_checksum <= x"ea";
					when x"50" => i_checksum <= x"b7";
					when x"51" => i_checksum <= x"b0";
					when x"52" => i_checksum <= x"b9";
					when x"53" => i_checksum <= x"be";
					when x"54" => i_checksum <= x"ab";
					when x"55" => i_checksum <= x"ac";
					when x"56" => i_checksum <= x"a5";
					when x"57" => i_checksum <= x"a2";
					when x"58" => i_checksum <= x"8f";
					when x"59" => i_checksum <= x"88";
					when x"5a" => i_checksum <= x"81";
					when x"5b" => i_checksum <= x"86";
					when x"5c" => i_checksum <= x"93";
					when x"5d" => i_checksum <= x"94";
					when x"5e" => i_checksum <= x"9d";
					when x"5f" => i_checksum <= x"9a";
					when x"60" => i_checksum <= x"27";
					when x"61" => i_checksum <= x"20";
					when x"62" => i_checksum <= x"29";
					when x"63" => i_checksum <= x"2e";
					when x"64" => i_checksum <= x"3b";
					when x"65" => i_checksum <= x"3c";
					when x"66" => i_checksum <= x"35";
					when x"67" => i_checksum <= x"32";
					when x"68" => i_checksum <= x"1f";
					when x"69" => i_checksum <= x"18";
					when x"6a" => i_checksum <= x"11";
					when x"6b" => i_checksum <= x"16";
					when x"6c" => i_checksum <= x"03";
					when x"6d" => i_checksum <= x"04";
					when x"6e" => i_checksum <= x"0d";
					when x"6f" => i_checksum <= x"0a";
					when x"70" => i_checksum <= x"57";
					when x"71" => i_checksum <= x"50";
					when x"72" => i_checksum <= x"59";
					when x"73" => i_checksum <= x"5e";
					when x"74" => i_checksum <= x"4b";
					when x"75" => i_checksum <= x"4c";
					when x"76" => i_checksum <= x"45";
					when x"77" => i_checksum <= x"42";
					when x"78" => i_checksum <= x"6f";
					when x"79" => i_checksum <= x"68";
					when x"7a" => i_checksum <= x"61";
					when x"7b" => i_checksum <= x"66";
					when x"7c" => i_checksum <= x"73";
					when x"7d" => i_checksum <= x"74";
					when x"7e" => i_checksum <= x"7d";
					when x"7f" => i_checksum <= x"7a";
					when x"80" => i_checksum <= x"89";
					when x"81" => i_checksum <= x"8e";
					when x"82" => i_checksum <= x"87";
					when x"83" => i_checksum <= x"80";
					when x"84" => i_checksum <= x"95";
					when x"85" => i_checksum <= x"92";
					when x"86" => i_checksum <= x"9b";
					when x"87" => i_checksum <= x"9c";
					when x"88" => i_checksum <= x"b1";
					when x"89" => i_checksum <= x"b6";
					when x"8a" => i_checksum <= x"bf";
					when x"8b" => i_checksum <= x"b8";
					when x"8c" => i_checksum <= x"ad";
					when x"8d" => i_checksum <= x"aa";
					when x"8e" => i_checksum <= x"a3";
					when x"8f" => i_checksum <= x"a4";
					when x"90" => i_checksum <= x"f9";
					when x"91" => i_checksum <= x"fe";
					when x"92" => i_checksum <= x"f7";
					when x"93" => i_checksum <= x"f0";
					when x"94" => i_checksum <= x"e5";
					when x"95" => i_checksum <= x"e2";
					when x"96" => i_checksum <= x"eb";
					when x"97" => i_checksum <= x"ec";
					when x"98" => i_checksum <= x"c1";
					when x"99" => i_checksum <= x"c6";
					when x"9a" => i_checksum <= x"cf";
					when x"9b" => i_checksum <= x"c8";
					when x"9c" => i_checksum <= x"dd";
					when x"9d" => i_checksum <= x"da";
					when x"9e" => i_checksum <= x"d3";
					when x"9f" => i_checksum <= x"d4";
					when x"a0" => i_checksum <= x"69";
					when x"a1" => i_checksum <= x"6e";
					when x"a2" => i_checksum <= x"67";
					when x"a3" => i_checksum <= x"60";
					when x"a4" => i_checksum <= x"75";
					when x"a5" => i_checksum <= x"72";
					when x"a6" => i_checksum <= x"7b";
					when x"a7" => i_checksum <= x"7c";
					when x"a8" => i_checksum <= x"51";
					when x"a9" => i_checksum <= x"56";
					when x"aa" => i_checksum <= x"5f";
					when x"ab" => i_checksum <= x"58";
					when x"ac" => i_checksum <= x"4d";
					when x"ad" => i_checksum <= x"4a";
					when x"ae" => i_checksum <= x"43";
					when x"af" => i_checksum <= x"44";
					when x"b0" => i_checksum <= x"19";
					when x"b1" => i_checksum <= x"1e";
					when x"b2" => i_checksum <= x"17";
					when x"b3" => i_checksum <= x"10";
					when x"b4" => i_checksum <= x"05";
					when x"b5" => i_checksum <= x"02";
					when x"b6" => i_checksum <= x"0b";
					when x"b7" => i_checksum <= x"0c";
					when x"b8" => i_checksum <= x"21";
					when x"b9" => i_checksum <= x"26";
					when x"ba" => i_checksum <= x"2f";
					when x"bb" => i_checksum <= x"28";
					when x"bc" => i_checksum <= x"3d";
					when x"bd" => i_checksum <= x"3a";
					when x"be" => i_checksum <= x"33";
					when x"bf" => i_checksum <= x"34";
					when x"c0" => i_checksum <= x"4e";
					when x"c1" => i_checksum <= x"49";
					when x"c2" => i_checksum <= x"40";
					when x"c3" => i_checksum <= x"47";
					when x"c4" => i_checksum <= x"52";
					when x"c5" => i_checksum <= x"55";
					when x"c6" => i_checksum <= x"5c";
					when x"c7" => i_checksum <= x"5b";
					when x"c8" => i_checksum <= x"76";
					when x"c9" => i_checksum <= x"71";
					when x"ca" => i_checksum <= x"78";
					when x"cb" => i_checksum <= x"7f";
					when x"cc" => i_checksum <= x"6a";
					when x"cd" => i_checksum <= x"6d";
					when x"ce" => i_checksum <= x"64";
					when x"cf" => i_checksum <= x"63";
					when x"d0" => i_checksum <= x"3e";
					when x"d1" => i_checksum <= x"39";
					when x"d2" => i_checksum <= x"30";
					when x"d3" => i_checksum <= x"37";
					when x"d4" => i_checksum <= x"22";
					when x"d5" => i_checksum <= x"25";
					when x"d6" => i_checksum <= x"2c";
					when x"d7" => i_checksum <= x"2b";
					when x"d8" => i_checksum <= x"06";
					when x"d9" => i_checksum <= x"01";
					when x"da" => i_checksum <= x"08";
					when x"db" => i_checksum <= x"0f";
					when x"dc" => i_checksum <= x"1a";
					when x"dd" => i_checksum <= x"1d";
					when x"de" => i_checksum <= x"14";
					when x"df" => i_checksum <= x"13";
					when x"e0" => i_checksum <= x"ae";
					when x"e1" => i_checksum <= x"a9";
					when x"e2" => i_checksum <= x"a0";
					when x"e3" => i_checksum <= x"a7";
					when x"e4" => i_checksum <= x"b2";
					when x"e5" => i_checksum <= x"b5";
					when x"e6" => i_checksum <= x"bc";
					when x"e7" => i_checksum <= x"bb";
					when x"e8" => i_checksum <= x"96";
					when x"e9" => i_checksum <= x"91";
					when x"ea" => i_checksum <= x"98";
					when x"eb" => i_checksum <= x"9f";
					when x"ec" => i_checksum <= x"8a";
					when x"ed" => i_checksum <= x"8d";
					when x"ee" => i_checksum <= x"84";
					when x"ef" => i_checksum <= x"83";
					when x"f0" => i_checksum <= x"de";
					when x"f1" => i_checksum <= x"d9";
					when x"f2" => i_checksum <= x"d0";
					when x"f3" => i_checksum <= x"d7";
					when x"f4" => i_checksum <= x"c2";
					when x"f5" => i_checksum <= x"c5";
					when x"f6" => i_checksum <= x"cc";
					when x"f7" => i_checksum <= x"cb";
					when x"f8" => i_checksum <= x"e6";
					when x"f9" => i_checksum <= x"e1";
					when x"fa" => i_checksum <= x"e8";
					when x"fb" => i_checksum <= x"ef";
					when x"fc" => i_checksum <= x"fa";
					when x"fd" => i_checksum <= x"fd";
					when x"fe" => i_checksum <= x"f4";
					when x"ff" => i_checksum <= x"f3";
					when others => null;
				end case;
			else
				if update = '1' then
					i_checksum <= i_checksum xor data;
					load_table <= '1';
				end if;
				checksum <= i_checksum;
			end if;
			if init = '1' then
				i_checksum <= (others => '0');
			end if;
		end if;
	end process;

end Behavior;
